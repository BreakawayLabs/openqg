netcdf ocn_basin_cdl {

dimensions:
	strlen = 64;
	nl = 3;
	nlm1 = 2;
	out = 7;

variables:
	char name(strlen);

	integer nx, ny;
	integer ndx, ndy;
	integer nx1, ny1;
	double hm, h(nl);

	char topog(strlen);

	double rho;

	integer use_oml;

	integer use_qg;
	double bcco;
	double delek;
	double ah2(nl), ah4(nl);
	double gp(nlm1);
	char qg_state(strlen);

	char ent_cpl(strlen);

	integer compute_covar;

	integer compute_avges;
	double dtav;
	char avg_out(strlen);

	integer compute_subsample;
	double dtsubsamp;
	char p_file(strlen);
	char t_file(strlen);
	integer nsk;
	integer outfl(out);

	integer check_valids;
	double dtvalid;
	double max_tau;
	double max_wt;
	double max_st;
	double max_p;
	double max_q;

	integer print_summary;
	double dtprint;

	integer area_avg;

	integer monitor_qg;
	char qg_mon_out(strlen);

	integer monitor_ml;
	char ml_mon_out(strlen);

	double dtdiag;	
data:
	name = "southern_ocean";

	nx = 288;
	ny = 36;
	ndx = 8;
	ndy = 8;
	nx1 = 1;
	ny1 = 37;
	hm = 100.0;
	h = 300.0,  1100.0, 2600.0;

	topog = "soctopog.26deg.10km.new.nc";

	rho = 1.0e3;

	use_oml = 0;

	use_qg = 1;
	bcco  = 5.0;
	delek = 2.0;
	ah2 = 0.0,    0.0,    0.0;
	ah4 = 3.0e10, 3.0e10, 3.0e10;
	gp  =     5.0e-2,  2.5e-2;
	qg_state = "zero";

	ent_cpl = "zero";

	compute_covar = 0;

	compute_avges = 0;
	dtav = 1.0;
	avg_out = "avges_ocn.nc";

	compute_subsample = 1;
	dtsubsamp = 15.0;
	p_file = "ocpo.nc";
	t_file = "ocsst.nc";
	nsk = 4;
	outfl = 1, 1, 1, 1, 1, 1, 1;

	check_valids = 1;
	dtvalid = 0.25;
	max_tau = 10.0e0;
	max_wt = 1.0e-3;
	max_st = 90.0e0;
	max_p = 1.0e4;
	max_q = 0.05e0;

	print_summary = 1;
	dtprint = 1.0;

	area_avg = 0;

	monitor_qg = 1;
	qg_mon_out = "qgo_mon.nc";

	monitor_ml = 1;
	ml_mon_out = "oml_mon.nc";

	dtdiag = 1.0;

}