netcdf windstress {

variables:
	integer coupled;
	double cdat;
	integer tau_udiff;
data:
	coupled = 1;
	cdat = 1.3e-3;
	tau_udiff = 0;
}