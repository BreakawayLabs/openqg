netcdf so_coupled_topog_glam {

dimensions:
	strlen = 64;
	oc_nl = 3;
	at_nl = 3;

variables:
	integer nxt, nyt;
	double dx, dy;
	double x0, y0;
	integer cyclic;
	double lat, x1;

	integer use_ocean;

	integer use_atmos;
data:
	nxt = 288;
	nyt = 108;
	dx = 80.0e3;
	dy = 80.0e3;
	x0 = 0.0;
	y0 = 0.0;

	cyclic = 1;
	lat = -55.0;
	x1 = 0.0;

	use_atmos = 0;

	use_ocean = 1;
}