netcdf atm_basin_cdl {

dimensions:
	strlen = 64;
	nl = 3;
	nlm1 = 2;
	out = 7;
	narea = 6;

variables:
	char name(strlen);

	integer nx, ny;
	integer ndx, ndy;
	integer nx1, ny1;
	double hm, h(nl);

	char topog(strlen);

	double rho;

	integer use_aml;
	integer flux_n, flux_s;
	double st2d, st4d, ahmd;
	double cp;
	double hmamin, hmadmp, xcexp;

	double T_abs(nl);
	double fsbar, fspamp;
	double zopt_m, zopt(nl);
	double gamma, xlamda;
	char aml_state(strlen);

	integer use_qg;
	double bcco;
	double delek;
	double ah2(nl), ah4(nl);
	double gp(nlm1);
	char qg_state(strlen);

	char sst_cpl(strlen);
	char p1_cpl(strlen);
	char eta_cpl(strlen);
	char ent_cpl(strlen);

	integer compute_covar;

	integer compute_avges;
	double dtav;
	char avg_out(strlen);

	integer compute_subsample;
	double dtsubsamp;
	char p_file(strlen);
	char t_file(strlen);
	integer nsk;
	integer outfl(out);

	integer check_valids;
	double dtvalid;
	double max_tau;
	double max_wt;
	double max_st;
	double max_p;
	double max_q;

	integer print_summary;
	double dtprint;

	integer area_avg;
	double xhi(narea);
	double xlo(narea);
	double yhi(narea);
	double ylo(narea);
	char area_filename(strlen);

	integer monitor_qg;
	char qg_mon_out(strlen);

	integer monitor_ml;
	char ml_mon_out(strlen);

	double dtdiag;
data:
	name = "dg_atmos";

	nx = 128;
	ny = 64;
	ndx = 1;
	ndy = 1;
	nx1 = 1;
	ny1 = 1;
	hm = 1000.0;
	h = 2000.0, 3000.0, 4000.0;
	
	topog = "flat";

	rho = 1.0;

	use_aml = 1;
	flux_n = 0;
	flux_s = 0;
	st2d = 5.0e4;
	st4d = 3.0e14;
	ahmd = 2.0e5;
	cp = 1.0e3;
	hmamin = 100.0;
	hmadmp = 0.15;
	xcexp = 1.0;
	T_abs = 330.0,  340.0,  350.0;
	fsbar = -210.0;
	fspamp = 80.0;
	zopt_m = 200.0;
	zopt = 3.0e4,  3.0e4,  4.0e4;
	gamma = 1.0e-2;
	xlamda = 35.0;
	aml_state = "rbal";

	use_qg = 1;
	bcco  = 1.0;
	delek = 0.0;
	ah2 = 0.0,    0.0,    0.0;
	ah4 = 2.0e13, 2.0e13, 2.0e13;
	gp  =       1.2,    0.4;
	qg_state = "rbal";

	sst_cpl = "coupled";
	p1_cpl = "coupled";
	eta_cpl = "coupled";
	ent_cpl = "coupled";

	compute_covar = 0;

	compute_avges = 0;
	dtav = 0.125;
	avg_out = "avges_atm.nc";

	compute_subsample = 1;
	dtsubsamp = 3.0;
	p_file = "atpa.nc";
	t_file = "atast.nc";
	nsk = 1;
	outfl = 1, 1, 1, 1, 1, 1, 1;

	check_valids = 1;
	dtvalid = 0.1;
	max_tau = 10.0e0;
	max_wt = 1.0;
	max_st = 90.0e0;
	max_p = 1.0e7;
	max_q = 0.05e0;

	print_summary = 1;
	dtprint = 1.0;

	area_avg = 1;
	xlo =    0.0e3,    0.0e3, 6000.0e3, 6000.0e3, 10000.0e3, 10000.0e3;
	xhi = 5000.0e3, 5000.0e3, 9000.0e3, 9000.0e3, 15000.0e3, 15000.0e3;
	ylo = 1440.0e3, 3840.0e3, 1400.0e3, 3840.0e3,  1400.0e3,  3840.0e3;
	yhi = 3840.0e3, 6240.0e3, 3840.0e3, 6240.0e3,  3840.0e3,  6240.0e3;
	area_filename = "atm_areas.nc";

	monitor_qg = 1;
	qg_mon_out = "qga_mon.nc";

	monitor_ml = 1;
	ml_mon_out = "aml_mon.nc";

	dtdiag = 1.0;
}