netcdf clock {

variables:
	double dta;
	double tini;
	double trun;
	integer nstr;
	double resday;

data:
	dta = 300.0;
	tini = 0.0;
	trun = 0.027397260;
	nstr = 3;
	resday = 365.0;
}
